module test (
	input clock
);

reg [3:0] array[4] = '{4'd1, 4'd2, 4'd3, 4'd4};

endmodule
module test;